// file ID_EX.v

module ID_EX(
	input wire [31:0] ID_RS,
	input wire [31:0] ID_RT,
	input wire [4:0] ID_RD,
	input wire clock,
	output reg [31:0] EX_RS,
	output reg [31:0] EX_RT,
	output reg [4:0] EX_RD);
	
	
	
	
endmodule
